`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:15:42 11/06/2017 
// Design Name: 
// Module Name:    DCT_2D 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
///////////////////////////////////////////////
module DCT_2D( 

//Inputs
I00, I01, I02, I03, I04, I05, I06, I07,
I10, I11, I12, I13, I14, I15, I16, I17,
I20, I21, I22, I23, I24, I25, I26, I27,
I30, I31, I32, I33, I34, I35, I36, I37,
I40, I41, I42, I43, I44, I45, I46, I47,
I50, I51, I52, I53, I54, I55, I56, I57,
I60, I61, I62, I63, I64, I65, I66, I67,
I70, I71, I72, I73, I74, I75, I76, I77, aclk,

//Outputs

O00, O01, O02, O03, O04, O05, O06, O07,
O10, O11, O12, O13, O14, O15, O16, O17,
O20, O21, O22, O23, O24, O25, O26, O27,
O30, O31, O32, O33, O34, O35, O36, O37,
O40, O41, O42, O43, O44, O45, O46, O47,
O50, O51, O52, O53, O54, O55, O56, O57,
O60, O61, O62, O63, O64, O65, O66, O67,
O70, O71, O72, O73, O74, O75, O76, O77
);


input [31:0] 
I00, I01, I02, I03, I04, I05, I06, I07,
I10, I11, I12, I13, I14, I15, I16, I17,
I20, I21, I22, I23, I24, I25, I26, I27,
I30, I31, I32, I33, I34, I35, I36, I37,
I40, I41, I42, I43, I44, I45, I46, I47,
I50, I51, I52, I53, I54, I55, I56, I57,
I60, I61, I62, I63, I64, I65, I66, I67,
I70, I71, I72, I73, I74, I75, I76, I77;

input aclk;

output wire [31:0] 
O00, O01, O02, O03, O04, O05, O06, O07,
O10, O11, O12, O13, O14, O15, O16, O17,
O20, O21, O22, O23, O24, O25, O26, O27,
O30, O31, O32, O33, O34, O35, O36, O37,
O40, O41, O42, O43, O44, O45, O46, O47,
O50, O51, O52, O53, O54, O55, O56, O57,
O60, O61, O62, O63, O64, O65, O66, O67,
O70, O71, O72, O73, O74, O75, O76, O77;



wire [31:0] 
TO00, TO01, TO02, TO03, TO04, TO05, TO06, TO07,
TO10, TO11, TO12, TO13, TO14, TO15, TO16, TO17,
TO20, TO21, TO22, TO23, TO24, TO25, TO26, TO27,
TO30, TO31, TO32, TO33, TO34, TO35, TO36, TO37,
TO40, TO41, TO42, TO43, TO44, TO45, TO46, TO47,
TO50, TO51, TO52, TO53, TO54, TO55, TO56, TO57,
TO60, TO61, TO62, TO63, TO64, TO65, TO66, TO67,
TO70, TO71, TO72, TO73, TO74, TO75, TO76, TO77;


DCT_1D   Stage1_0(I00, I01, I02, I03, I04, I05, I06, I07, TO00, TO01, TO02, TO03, TO04, TO05, TO06, TO07, aclk);
DCT_1D   Stage1_1(I10, I11, I12, I13, I14, I15, I16, I17, TO10, TO11, TO12, TO13, TO14, TO15, TO16, TO17, aclk);
DCT_1D   Stage1_2(I20, I21, I22, I23, I24, I25, I26, I27, TO20, TO21, TO22, TO23, TO24, TO25, TO26, TO27, aclk);
DCT_1D   Stage1_3(I30, I31, I32, I33, I34, I35, I36, I37, TO30, TO31, TO32, TO33, TO34, TO35, TO36, TO37, aclk);
DCT_1D   Stage1_4(I40, I41, I42, I43, I44, I45, I46, I47, TO40, TO41, TO42, TO43, TO44, TO45, TO46, TO47, aclk);
DCT_1D   Stage1_5(I50, I51, I52, I53, I54, I55, I56, I57, TO50, TO51, TO52, TO53, TO54, TO55, TO56, TO57, aclk);
DCT_1D   Stage1_6(I60, I61, I62, I63, I64, I65, I66, I67, TO60, TO61, TO62, TO63, TO64, TO65, TO66, TO67, aclk);
DCT_1D   Stage1_7(I70, I71, I72, I73, I74, I75, I76, I77, TO70, TO71, TO72, TO73, TO74, TO75, TO76, TO77, aclk);


DCT_1D   Stage2_0(TO00, TO10, TO20, TO30, TO40, TO50, TO60, TO70, O00, O01, O02, O03, O04, O05, O06,  O07, aclk);
DCT_1D   Stage2_1(TO01, TO11, TO21, TO31, TO41, TO51, TO61, TO71, O10, O11, O12, O13, O14, O15, O16,  O17, aclk);
DCT_1D   Stage2_2(TO02, TO12, TO22, TO32, TO42, TO52, TO62, TO72, O20, O21, O22, O23, O24, O25, O26,  O27, aclk);
DCT_1D   Stage2_3(TO03, TO13, TO23, TO33, TO43, TO53, TO63, TO73, O30, O31, O32, O33, O34, O35, O36,  O37, aclk);
DCT_1D   Stage2_4(TO04, TO14, TO24, TO34, TO44, TO54, TO64, TO74, O40, O41, O42, O43, O44, O45, O46,  O47, aclk);
DCT_1D   Stage2_5(TO05, TO15, TO25, TO35, TO45, TO55, TO65, TO75, O50, O51, O52, O53, O54, O55, O56,  O57, aclk);
DCT_1D   Stage2_6(TO06, TO16, TO26, TO36, TO46, TO56, TO66, TO76, O60, O61, O62, O63, O64, O65, O66,  O67, aclk);
DCT_1D   Stage2_7(TO07, TO17, TO27, TO37, TO47, TO57, TO67, TO77, O70, O71, O72, O73, O74, O75, O76,  O77, aclk);



//-----------QUANTIZATION--------------------------//


endmodule

